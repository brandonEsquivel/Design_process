* First line is ignored

*** SUBCIRCUIT NAND3 FROM CELL NAND3{lay}
.SUBCKT NAND3 A B C gnd vdd Y_NAND3
Mnmos@4 net@17 A gnd gnd N L=0.4U W=1U
Mnmos@5 net@16 B net@17 gnd N L=0.4U W=1U
Mnmos@6 Y_NAND3 C net@16 gnd N L=0.4U W=1U
Mpmos@3 Y_NAND3 A vdd vdd P L=0.4U W=2U
Mpmos@4 vdd B Y_NAND3 vdd P L=0.4U W=2U
Mpmos@5 Y_NAND3 C vdd vdd P L=0.4U W=2U
.ENDS NAND3
