module counter ( gnd, vdd, ENABLE, RESET, clk, D, MODO, Q, RCO, LOAD);

input gnd, vdd;
input ENABLE;
input RESET;
input clk;
output RCO;
input [31:0] D;
input [1:0] MODO;
output [31:0] Q;
output [7:0] LOAD;

	BUFX4 BUFX4_1 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf8) );
	BUFX4 BUFX4_2 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf7) );
	BUFX4 BUFX4_3 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf6) );
	BUFX4 BUFX4_4 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf5) );
	BUFX4 BUFX4_5 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf4) );
	BUFX4 BUFX4_6 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf3) );
	BUFX4 BUFX4_7 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf2) );
	BUFX4 BUFX4_8 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf1) );
	BUFX4 BUFX4_9 ( .gnd(gnd), .vdd(vdd), .A(clk), .Y(clk_bF_buf0) );
	BUFX4 BUFX4_10 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf7) );
	BUFX4 BUFX4_11 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf6) );
	BUFX4 BUFX4_12 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf5) );
	BUFX4 BUFX4_13 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf4) );
	BUFX4 BUFX4_14 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf3) );
	BUFX4 BUFX4_15 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf2) );
	BUFX4 BUFX4_16 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf1) );
	BUFX4 BUFX4_17 ( .gnd(gnd), .vdd(vdd), .A(RESET), .Y(RESET_bF_buf0) );
	NAND2X1 NAND2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_361_), .Y(_369_) );
	NAND2X1 NAND2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_396_), .Y(_370_) );
	AOI22X1 AOI22X1_1 ( .gnd(gnd), .vdd(vdd), .A(D_reg_23_), .B(_331_), .C(_370_), .D(_338_), .Y(_371_) );
	AOI21X1 AOI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_371_), .B(_386_), .C(_328_), .Y(_325__3_) );
	DFFPOSX1 DFFPOSX1_1 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_325__0_), .Q(_82__24_) );
	DFFPOSX1 DFFPOSX1_2 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_355__1_), .Q(_82__25_) );
	DFFPOSX1 DFFPOSX1_3 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_355__2_), .Q(_82__26_) );
	DFFPOSX1 DFFPOSX1_4 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_355__3_), .Q(_82__27_) );
	DFFPOSX1 DFFPOSX1_5 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_326_), .Q(cont4b_5_RCO) );
	DFFPOSX1 DFFPOSX1_6 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_324_), .Q(cont4b_5_LOAD) );
	INVX1 INVX1_1 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .Y(_375_) );
	NAND2X1 NAND2X1_3 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_402_), .Y(_376_) );
	INVX1 INVX1_2 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_6__0_), .Y(_377_) );
	INVX1 INVX1_3 ( .gnd(gnd), .vdd(vdd), .A(_406_), .Y(_378_) );
	NOR2X1 NOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_405_), .Y(_379_) );
	INVX1 INVX1_4 ( .gnd(gnd), .vdd(vdd), .A(_408_), .Y(_380_) );
	NOR2X1 NOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_403_), .B(_407_), .Y(_372_) );
	NOR2X1 NOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_7__1_), .B(_404_), .Y(_381_) );
	AOI21X1 AOI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_390_), .B(_392_), .C(_358_), .Y(_382_) );
	INVX1 INVX1_5 ( .gnd(gnd), .vdd(vdd), .A(_382_), .Y(_383_) );
	NOR2X1 NOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_82__27_), .B(_383_), .Y(_384_) );
	NAND2X1 NAND2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .B(_82__29_), .Y(_385_) );
	NOR2X1 NOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_7__0_), .B(_405_), .Y(_386_) );
	INVX1 INVX1_6 ( .gnd(gnd), .vdd(vdd), .A(_82__27_), .Y(_387_) );
	INVX1 INVX1_7 ( .gnd(gnd), .vdd(vdd), .A(_416_), .Y(_388_) );
	NOR2X1 NOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_82__31_), .B(_417_), .Y(_389_) );
	NAND3X1 NAND3X1_1 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_388_), .C(_389_), .Y(_390_) );
	INVX1 INVX1_8 ( .gnd(gnd), .vdd(vdd), .A(_82__28_), .Y(_391_) );
	NOR2X1 NOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_7__0_), .B(MODO_reg_7__1_), .Y(_392_) );
	AND2X2 AND2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_82__31_), .Y(_393_) );
	NAND2X1 NAND2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_82__26_), .B(_406_), .Y(_394_) );
	NOR2X1 NOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_82__28_), .B(_421_), .Y(_395_) );
	AOI22X1 AOI22X1_2 ( .gnd(gnd), .vdd(vdd), .A(_393_), .B(_361_), .C(_363_), .D(_391_), .Y(_396_) );
	AOI21X1 AOI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_395_), .C(_358_), .Y(_374_) );
	NAND2X1 NAND2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_82__29_), .B(_82__28_), .Y(_397_) );
	INVX1 INVX1_9 ( .gnd(gnd), .vdd(vdd), .A(_82__24_), .Y(_398_) );
	OAI21X1 OAI21X1_1 ( .gnd(gnd), .vdd(vdd), .A(_377_), .B(_378_), .C(_388_), .Y(_399_) );
	AOI21X1 AOI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_82__29_), .B(_82__28_), .C(_82__30_), .Y(_373__0_) );
	INVX1 INVX1_10 ( .gnd(gnd), .vdd(vdd), .A(_82__25_), .Y(_400_) );
	NOR2X1 NOR2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .Y(_401_) );
	NOR2X1 NOR2X1_10 ( .gnd(gnd), .vdd(vdd), .A(_88_), .B(_92_), .Y(_402_) );
	NAND2X1 NAND2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_428_), .B(_427_), .Y(_403_) );
	OR2X2 OR2X2_1 ( .gnd(gnd), .vdd(vdd), .A(_409_), .B(_413_), .Y(_404_) );
	AOI22X1 AOI22X1_3 ( .gnd(gnd), .vdd(vdd), .A(_394_), .B(_374_), .C(_404_), .D(_393_), .Y(_405_) );
	AOI21X1 AOI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(_423_), .B(_414_), .C(_403_), .Y(_373__1_) );
	OAI21X1 OAI21X1_2 ( .gnd(gnd), .vdd(vdd), .A(_398_), .B(_388_), .C(_389_), .Y(_406_) );
	OAI21X1 OAI21X1_3 ( .gnd(gnd), .vdd(vdd), .A(_82__26_), .B(_378_), .C(_82__27_), .Y(_407_) );
	OAI21X1 OAI21X1_4 ( .gnd(gnd), .vdd(vdd), .A(_404_), .B(_405_), .C(_425_), .Y(_408_) );
	NAND3X1 NAND3X1_2 ( .gnd(gnd), .vdd(vdd), .A(_410_), .B(_411_), .C(_412_), .Y(_409_) );
	OAI21X1 OAI21X1_5 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_7__0_), .B(_405_), .C(_433_), .Y(_410_) );
	NAND2X1 NAND2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_417_), .Y(_411_) );
	AOI22X1 AOI22X1_4 ( .gnd(gnd), .vdd(vdd), .A(D_reg_26_), .B(_361_), .C(_363_), .D(_397_), .Y(_412_) );
	AOI21X1 AOI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_424_), .B(_426_), .C(_403_), .Y(_373__2_) );
	XOR2X1 XOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_382_), .B(_82__27_), .Y(_413_) );
	NAND3X1 NAND3X1_3 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .B(_82__29_), .C(_82__28_), .Y(_414_) );
	XNOR2X1 XNOR2X1_1 ( .gnd(gnd), .vdd(vdd), .A(_414_), .B(_82__27_), .Y(_415_) );
	AOI22X1 AOI22X1_5 ( .gnd(gnd), .vdd(vdd), .A(_420_), .B(_422_), .C(_415_), .D(_418_), .Y(_416_) );
	NAND2X1 NAND2X1_9 ( .gnd(gnd), .vdd(vdd), .A(_413_), .B(_441_), .Y(_417_) );
	NAND2X1 NAND2X1_10 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(_417_), .Y(_418_) );
	AOI22X1 AOI22X1_6 ( .gnd(gnd), .vdd(vdd), .A(D_reg_27_), .B(_406_), .C(_408_), .D(_429_), .Y(_419_) );
	AOI21X1 AOI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_431_), .C(_403_), .Y(_373__3_) );
	DFFPOSX1 DFFPOSX1_7 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_400__0_), .Q(_82__28_) );
	DFFPOSX1 DFFPOSX1_8 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_400__1_), .Q(_82__29_) );
	DFFPOSX1 DFFPOSX1_9 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_400__2_), .Q(_82__30_) );
	DFFPOSX1 DFFPOSX1_10 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_400__3_), .Q(_82__31_) );
	DFFPOSX1 DFFPOSX1_11 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_401_), .Q(cont4b_6_RCO) );
	DFFPOSX1 DFFPOSX1_12 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_399_), .Q(cont4b_6_LOAD) );
	INVX1 INVX1_11 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .Y(_423_) );
	NAND2X1 NAND2X1_11 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(_423_), .Y(_424_) );
	INVX1 INVX1_12 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_7__0_), .Y(_425_) );
	INVX1 INVX1_13 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_7__1_), .Y(_426_) );
	NOR2X1 NOR2X1_11 ( .gnd(gnd), .vdd(vdd), .A(MODO[1]), .B(_89_), .Y(_427_) );
	INVX1 INVX1_14 ( .gnd(gnd), .vdd(vdd), .A(_427_), .Y(_428_) );
	NOR2X1 NOR2X1_12 ( .gnd(gnd), .vdd(vdd), .A(_82__1_), .B(_82__0_), .Y(_420_) );
	NOR2X1 NOR2X1_13 ( .gnd(gnd), .vdd(vdd), .A(MODO[0]), .B(_90_), .Y(_429_) );
	AOI21X1 AOI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_437_), .C(_403_), .Y(_430_) );
	INVX1 INVX1_15 ( .gnd(gnd), .vdd(vdd), .A(_430_), .Y(_431_) );
	NOR2X1 NOR2X1_14 ( .gnd(gnd), .vdd(vdd), .A(_82__3_), .B(_102_), .Y(_432_) );
	NAND2X1 NAND2X1_12 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(_432_), .Y(_433_) );
	NOR2X1 NOR2X1_15 ( .gnd(gnd), .vdd(vdd), .A(MODO[0]), .B(MODO[1]), .Y(_434_) );
	INVX1 INVX1_16 ( .gnd(gnd), .vdd(vdd), .A(_82__31_), .Y(_435_) );
	INVX1 INVX1_17 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .Y(_436_) );
	NOR2X1 NOR2X1_16 ( .gnd(gnd), .vdd(vdd), .A(_82__0_), .B(_106_), .Y(_437_) );
	NAND3X1 NAND3X1_4 ( .gnd(gnd), .vdd(vdd), .A(_435_), .B(_15_), .C(_16_), .Y(_438_) );
	INVX1 INVX1_18 ( .gnd(gnd), .vdd(vdd), .A(_438_), .Y(_439_) );
	NOR2X1 NOR2X1_17 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .Y(_440_) );
	AND2X2 AND2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_82__3_), .Y(_441_) );
	NAND2X1 NAND2X1_13 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(_82__29_), .Y(_442_) );
	NOR2X1 NOR2X1_18 ( .gnd(gnd), .vdd(vdd), .A(_133_), .B(_137_), .Y(_443_) );
	AOI22X1 AOI22X1_7 ( .gnd(gnd), .vdd(vdd), .A(_441_), .B(_406_), .C(_408_), .D(_436_), .Y(_444_) );
	AOI21X1 AOI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(_443_), .B(_440_), .C(_403_), .Y(_422_) );
	NAND2X1 NAND2X1_14 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(_427_), .Y(_445_) );
	INVX1 INVX1_19 ( .gnd(gnd), .vdd(vdd), .A(_82__28_), .Y(_446_) );
	OAI21X1 OAI21X1_6 ( .gnd(gnd), .vdd(vdd), .A(_419_), .B(_433_), .C(_434_), .Y(_447_) );
	AOI21X1 AOI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(_82__1_), .B(_82__0_), .C(_82__2_), .Y(_421__0_) );
	INVX1 INVX1_20 ( .gnd(gnd), .vdd(vdd), .A(_82__29_), .Y(_448_) );
	NOR2X1 NOR2X1_19 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_1__1_), .B(_134_), .Y(_449_) );
	NOR2X1 NOR2X1_20 ( .gnd(gnd), .vdd(vdd), .A(_82__5_), .B(_82__4_), .Y(_450_) );
	NAND2X1 NAND2X1_15 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(_450_), .Y(_451_) );
	OR2X2 OR2X2_2 ( .gnd(gnd), .vdd(vdd), .A(_82__29_), .B(_82__28_), .Y(_452_) );
	AOI22X1 AOI22X1_8 ( .gnd(gnd), .vdd(vdd), .A(_439_), .B(_419_), .C(_415_), .D(_438_), .Y(_453_) );
	AOI21X1 AOI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(_108_), .B(_99_), .C(_88_), .Y(_421__1_) );
	OAI21X1 OAI21X1_7 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .B(_427_), .C(_82__31_), .Y(_454_) );
	OAI21X1 OAI21X1_8 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_18_), .C(_19_), .Y(_455_) );
	OAI21X1 OAI21X1_9 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_20_), .C(_21_), .Y(_456_) );
	NAND3X1 NAND3X1_5 ( .gnd(gnd), .vdd(vdd), .A(cont4b_3_RCO), .B(_15_), .C(_17_), .Y(_457_) );
	OAI21X1 OAI21X1_10 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_22_), .C(_23_), .Y(_458_) );
	NAND2X1 NAND2X1_16 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(_457_), .Y(_459_) );
	AOI22X1 AOI22X1_9 ( .gnd(gnd), .vdd(vdd), .A(D_reg_30_), .B(_406_), .C(_408_), .D(_442_), .Y(_460_) );
	AOI21X1 AOI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(_109_), .B(_111_), .C(_88_), .Y(_421__2_) );
	XOR2X1 XOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_430_), .B(_82__31_), .Y(_461_) );
	NAND3X1 NAND3X1_6 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .B(_15_), .C(_16_), .Y(_462_) );
	XNOR2X1 XNOR2X1_2 ( .gnd(gnd), .vdd(vdd), .A(_462_), .B(_82__31_), .Y(_463_) );
	AOI22X1 AOI22X1_10 ( .gnd(gnd), .vdd(vdd), .A(_105_), .B(_107_), .C(_100_), .D(_103_), .Y(_464_) );
	NAND2X1 NAND2X1_17 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(_457_), .Y(_465_) );
	NAND2X1 NAND2X1_18 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(_465_), .Y(_466_) );
	AOI22X1 AOI22X1_11 ( .gnd(gnd), .vdd(vdd), .A(D_reg_1_), .B(_91_), .C(_93_), .D(_114_), .Y(_467_) );
	AOI21X1 AOI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(_115_), .B(_116_), .C(_88_), .Y(_421__3_) );
	DFFPOSX1 DFFPOSX1_13 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_7_), .Q(_82__28_) );
	DFFPOSX1 DFFPOSX1_14 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_8_), .Q(_82__29_) );
	DFFPOSX1 DFFPOSX1_15 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_1_), .Q(_82__30_) );
	DFFPOSX1 DFFPOSX1_16 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_2_), .Q(_82__31_) );
	DFFPOSX1 DFFPOSX1_17 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_9_), .Q(_83_) );
	DFFPOSX1 DFFPOSX1_18 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_10_), .Q(cont4b_7_LOAD) );
	INVX4 INVX4_1 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .Y(_15_) );
	INVX2 INVX2_1 ( .gnd(gnd), .vdd(vdd), .A(MODO[0]), .Y(_16_) );
	NAND3X1 NAND3X1_7 ( .gnd(gnd), .vdd(vdd), .A(cont4b_1_RCO), .B(_15_), .C(_17_), .Y(_11_) );
	INVX2 INVX2_2 ( .gnd(gnd), .vdd(vdd), .A(MODO[1]), .Y(_17_) );
	NAND3X1 NAND3X1_8 ( .gnd(gnd), .vdd(vdd), .A(cont4b_3_RCO), .B(_15_), .C(_16_), .Y(_13_) );
	NAND3X1 NAND3X1_9 ( .gnd(gnd), .vdd(vdd), .A(cont4b_2_RCO), .B(_15_), .C(_17_), .Y(_1_) );
	NAND3X1 NAND3X1_10 ( .gnd(gnd), .vdd(vdd), .A(cont4b_6_RCO), .B(_15_), .C(_16_), .Y(_2_) );
	NAND3X1 NAND3X1_11 ( .gnd(gnd), .vdd(vdd), .A(cont4b_6_RCO), .B(_15_), .C(_17_), .Y(_9_) );
	NAND3X1 NAND3X1_12 ( .gnd(gnd), .vdd(vdd), .A(cont4b_2_RCO), .B(_15_), .C(_16_), .Y(_10_) );
	NAND3X1 NAND3X1_13 ( .gnd(gnd), .vdd(vdd), .A(cont4b_5_RCO), .B(_15_), .C(_17_), .Y(_12_) );
	NAND3X1 NAND3X1_14 ( .gnd(gnd), .vdd(vdd), .A(cont4b_6_RCO), .B(_15_), .C(_16_), .Y(_14_) );
	INVX1 INVX1_21 ( .gnd(gnd), .vdd(vdd), .A(_82__0_), .Y(_18_) );
	NAND2X1 NAND2X1_19 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(D[0]), .Y(_19_) );
	OAI21X1 OAI21X1_11 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_24_), .C(_25_), .Y(_0__0_) );
	INVX1 INVX1_22 ( .gnd(gnd), .vdd(vdd), .A(_82__1_), .Y(_20_) );
	NAND2X1 NAND2X1_20 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(D[1]), .Y(_21_) );
	OAI21X1 OAI21X1_12 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_26_), .C(_27_), .Y(_0__1_) );
	INVX1 INVX1_23 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .Y(_22_) );
	NAND2X1 NAND2X1_21 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(D[2]), .Y(_23_) );
	OAI21X1 OAI21X1_13 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_28_), .C(_29_), .Y(_0__2_) );
	INVX1 INVX1_24 ( .gnd(gnd), .vdd(vdd), .A(_82__3_), .Y(_24_) );
	NAND2X1 NAND2X1_22 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(D[3]), .Y(_25_) );
	OAI21X1 OAI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_30_), .C(_31_), .Y(_0__3_) );
	INVX1 INVX1_25 ( .gnd(gnd), .vdd(vdd), .A(_82__4_), .Y(_26_) );
	NAND2X1 NAND2X1_23 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(D[4]), .Y(_27_) );
	OAI21X1 OAI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_32_), .C(_33_), .Y(_0__4_) );
	INVX1 INVX1_26 ( .gnd(gnd), .vdd(vdd), .A(_82__5_), .Y(_28_) );
	NAND2X1 NAND2X1_24 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(D[5]), .Y(_29_) );
	OAI21X1 OAI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_34_), .C(_35_), .Y(_0__5_) );
	INVX1 INVX1_27 ( .gnd(gnd), .vdd(vdd), .A(_82__6_), .Y(_30_) );
	NAND2X1 NAND2X1_25 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(D[6]), .Y(_31_) );
	OAI21X1 OAI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_36_), .C(_37_), .Y(_0__6_) );
	INVX1 INVX1_28 ( .gnd(gnd), .vdd(vdd), .A(_82__7_), .Y(_32_) );
	NAND2X1 NAND2X1_26 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(D[7]), .Y(_33_) );
	OAI21X1 OAI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_38_), .C(_39_), .Y(_0__7_) );
	INVX1 INVX1_29 ( .gnd(gnd), .vdd(vdd), .A(_82__8_), .Y(_34_) );
	NAND2X1 NAND2X1_27 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(D[8]), .Y(_35_) );
	OAI21X1 OAI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_40_), .C(_41_), .Y(_0__8_) );
	INVX1 INVX1_30 ( .gnd(gnd), .vdd(vdd), .A(_82__9_), .Y(_36_) );
	NAND2X1 NAND2X1_28 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(D[9]), .Y(_37_) );
	OAI21X1 OAI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_42_), .C(_43_), .Y(_0__9_) );
	INVX1 INVX1_31 ( .gnd(gnd), .vdd(vdd), .A(_82__10_), .Y(_38_) );
	NAND2X1 NAND2X1_29 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(D[10]), .Y(_39_) );
	OAI21X1 OAI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_44_), .C(_45_), .Y(_0__10_) );
	INVX1 INVX1_32 ( .gnd(gnd), .vdd(vdd), .A(_82__11_), .Y(_40_) );
	NAND2X1 NAND2X1_30 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(D[11]), .Y(_41_) );
	OAI21X1 OAI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_46_), .C(_47_), .Y(_0__11_) );
	INVX1 INVX1_33 ( .gnd(gnd), .vdd(vdd), .A(_82__24_), .Y(_42_) );
	NAND2X1 NAND2X1_31 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(D[12]), .Y(_43_) );
	OAI21X1 OAI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_48_), .C(_49_), .Y(_0__12_) );
	INVX1 INVX1_34 ( .gnd(gnd), .vdd(vdd), .A(_82__25_), .Y(_44_) );
	NAND2X1 NAND2X1_32 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(D[13]), .Y(_45_) );
	OAI21X1 OAI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_50_), .C(_51_), .Y(_0__13_) );
	INVX1 INVX1_35 ( .gnd(gnd), .vdd(vdd), .A(_82__26_), .Y(_46_) );
	NAND2X1 NAND2X1_33 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(D[14]), .Y(_47_) );
	OAI21X1 OAI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_52_), .C(_53_), .Y(_0__14_) );
	INVX1 INVX1_36 ( .gnd(gnd), .vdd(vdd), .A(_82__27_), .Y(_48_) );
	NAND2X1 NAND2X1_34 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(D[15]), .Y(_49_) );
	OAI21X1 OAI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_54_), .C(_55_), .Y(_0__15_) );
	INVX1 INVX1_37 ( .gnd(gnd), .vdd(vdd), .A(_82__28_), .Y(_50_) );
	NAND2X1 NAND2X1_35 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(D[16]), .Y(_51_) );
	OAI21X1 OAI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_56_), .C(_57_), .Y(_0__16_) );
	INVX1 INVX1_38 ( .gnd(gnd), .vdd(vdd), .A(_82__29_), .Y(_52_) );
	NAND2X1 NAND2X1_36 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(D[17]), .Y(_53_) );
	OAI21X1 OAI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_58_), .C(_59_), .Y(_0__17_) );
	INVX1 INVX1_39 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .Y(_54_) );
	NAND2X1 NAND2X1_37 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(D[18]), .Y(_55_) );
	OAI21X1 OAI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_60_), .C(_61_), .Y(_0__18_) );
	INVX1 INVX1_40 ( .gnd(gnd), .vdd(vdd), .A(_82__31_), .Y(_56_) );
	NAND2X1 NAND2X1_38 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .B(D[19]), .Y(_57_) );
	OAI21X1 OAI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_62_), .C(_63_), .Y(_0__19_) );
	INVX1 INVX1_41 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf5), .Y(_58_) );
	NAND2X1 NAND2X1_39 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .B(D[20]), .Y(_59_) );
	OAI21X1 OAI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_64_), .C(_65_), .Y(_0__20_) );
	INVX1 INVX1_42 ( .gnd(gnd), .vdd(vdd), .A(MODO[0]), .Y(_60_) );
	NAND2X1 NAND2X1_40 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .B(D[21]), .Y(_61_) );
	OAI21X1 OAI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_66_), .C(_67_), .Y(_0__21_) );
	INVX1 INVX1_43 ( .gnd(gnd), .vdd(vdd), .A(_91_), .Y(_62_) );
	NAND2X1 NAND2X1_41 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .B(D[22]), .Y(_63_) );
	OAI21X1 OAI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_68_), .C(_69_), .Y(_0__22_) );
	INVX1 INVX1_44 ( .gnd(gnd), .vdd(vdd), .A(_93_), .Y(_64_) );
	NAND2X1 NAND2X1_42 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_87_), .Y(_65_) );
	OAI21X1 OAI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_70_), .C(_71_), .Y(_0__23_) );
	INVX1 INVX1_45 ( .gnd(gnd), .vdd(vdd), .A(_82__3_), .Y(_66_) );
	NAND2X1 NAND2X1_43 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .B(_82__1_), .Y(_67_) );
	OAI21X1 OAI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_72_), .C(_73_), .Y(_0__24_) );
	INVX1 INVX1_46 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .Y(_68_) );
	NAND2X1 NAND2X1_44 ( .gnd(gnd), .vdd(vdd), .A(D_reg_0_), .B(_91_), .Y(_69_) );
	OAI21X1 OAI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .B(_74_), .C(_75_), .Y(_0__25_) );
	INVX1 INVX1_47 ( .gnd(gnd), .vdd(vdd), .A(_101_), .Y(_70_) );
	NAND2X1 NAND2X1_45 ( .gnd(gnd), .vdd(vdd), .A(_82__1_), .B(_82__0_), .Y(_71_) );
	OAI21X1 OAI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .B(_76_), .C(_77_), .Y(_0__26_) );
	INVX1 INVX1_48 ( .gnd(gnd), .vdd(vdd), .A(_82__0_), .Y(_72_) );
	NAND2X1 NAND2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_113_), .B(_112_), .Y(_73_) );
	OAI21X1 OAI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .B(_78_), .C(_79_), .Y(_0__27_) );
	INVX1 INVX1_49 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf4), .Y(_74_) );
	NAND2X1 NAND2X1_47 ( .gnd(gnd), .vdd(vdd), .A(_117_), .B(_102_), .Y(_75_) );
	OAI21X1 OAI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf6), .B(_80_), .C(_81_), .Y(_0__28_) );
	INVX1 INVX1_50 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_1__0_), .Y(_76_) );
	NAND2X1 NAND2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_98_), .B(_126_), .Y(_77_) );
	OAI21X1 OAI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_89_), .B(_90_), .C(_110_), .Y(_0__29_) );
	INVX1 INVX1_51 ( .gnd(gnd), .vdd(vdd), .A(_136_), .Y(_78_) );
	NAND2X1 NAND2X1_49 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_132_), .Y(_79_) );
	OAI21X1 OAI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(MODO[0]), .B(_90_), .C(_118_), .Y(_0__30_) );
	INVX1 INVX1_52 ( .gnd(gnd), .vdd(vdd), .A(_138_), .Y(_80_) );
	NAND2X1 NAND2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_82__6_), .B(_82__5_), .Y(_81_) );
	OAI21X1 OAI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_104_), .B(_118_), .C(_119_), .Y(_0__31_) );
	NAND3X1 NAND3X1_15 ( .gnd(gnd), .vdd(vdd), .A(cont4b_0_RCO), .B(_15_), .C(_17_), .Y(_3_) );
	NAND3X1 NAND3X1_16 ( .gnd(gnd), .vdd(vdd), .A(cont4b_5_RCO), .B(_15_), .C(_16_), .Y(_4_) );
	NAND3X1 NAND3X1_17 ( .gnd(gnd), .vdd(vdd), .A(cont4b_4_RCO), .B(_15_), .C(_17_), .Y(_5_) );
	NAND3X1 NAND3X1_18 ( .gnd(gnd), .vdd(vdd), .A(_95_), .B(_96_), .C(_97_), .Y(_6_) );
	NAND3X1 NAND3X1_19 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .B(_82__1_), .C(_82__0_), .Y(_7_) );
	NAND3X1 NAND3X1_20 ( .gnd(gnd), .vdd(vdd), .A(_140_), .B(_141_), .C(_142_), .Y(_8_) );
	BUFX2 BUFX2_1 ( .gnd(gnd), .vdd(vdd), .A(cont4b_0_LOAD), .Y(LOAD[0]) );
	BUFX2 BUFX2_2 ( .gnd(gnd), .vdd(vdd), .A(cont4b_1_LOAD), .Y(LOAD[1]) );
	BUFX2 BUFX2_3 ( .gnd(gnd), .vdd(vdd), .A(cont4b_2_LOAD), .Y(LOAD[2]) );
	BUFX2 BUFX2_4 ( .gnd(gnd), .vdd(vdd), .A(cont4b_3_LOAD), .Y(LOAD[3]) );
	BUFX2 BUFX2_5 ( .gnd(gnd), .vdd(vdd), .A(cont4b_4_LOAD), .Y(LOAD[4]) );
	BUFX2 BUFX2_6 ( .gnd(gnd), .vdd(vdd), .A(cont4b_5_LOAD), .Y(LOAD[5]) );
	BUFX2 BUFX2_7 ( .gnd(gnd), .vdd(vdd), .A(cont4b_6_LOAD), .Y(LOAD[6]) );
	BUFX2 BUFX2_8 ( .gnd(gnd), .vdd(vdd), .A(cont4b_7_LOAD), .Y(LOAD[7]) );
	BUFX2 BUFX2_9 ( .gnd(gnd), .vdd(vdd), .A(_82__0_), .Y(Q[0]) );
	BUFX2 BUFX2_10 ( .gnd(gnd), .vdd(vdd), .A(_82__1_), .Y(Q[1]) );
	BUFX2 BUFX2_11 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .Y(Q[2]) );
	BUFX2 BUFX2_12 ( .gnd(gnd), .vdd(vdd), .A(_82__3_), .Y(Q[3]) );
	BUFX2 BUFX2_13 ( .gnd(gnd), .vdd(vdd), .A(_82__4_), .Y(Q[4]) );
	BUFX2 BUFX2_14 ( .gnd(gnd), .vdd(vdd), .A(_82__5_), .Y(Q[5]) );
	BUFX2 BUFX2_15 ( .gnd(gnd), .vdd(vdd), .A(_82__6_), .Y(Q[6]) );
	BUFX2 BUFX2_16 ( .gnd(gnd), .vdd(vdd), .A(_82__7_), .Y(Q[7]) );
	BUFX2 BUFX2_17 ( .gnd(gnd), .vdd(vdd), .A(_82__8_), .Y(Q[8]) );
	BUFX2 BUFX2_18 ( .gnd(gnd), .vdd(vdd), .A(_82__9_), .Y(Q[9]) );
	BUFX2 BUFX2_19 ( .gnd(gnd), .vdd(vdd), .A(_82__10_), .Y(Q[10]) );
	BUFX2 BUFX2_20 ( .gnd(gnd), .vdd(vdd), .A(_82__11_), .Y(Q[11]) );
	BUFX2 BUFX2_21 ( .gnd(gnd), .vdd(vdd), .A(_82__12_), .Y(Q[12]) );
	BUFX2 BUFX2_22 ( .gnd(gnd), .vdd(vdd), .A(_82__13_), .Y(Q[13]) );
	BUFX2 BUFX2_23 ( .gnd(gnd), .vdd(vdd), .A(_82__14_), .Y(Q[14]) );
	BUFX2 BUFX2_24 ( .gnd(gnd), .vdd(vdd), .A(_82__15_), .Y(Q[15]) );
	BUFX2 BUFX2_25 ( .gnd(gnd), .vdd(vdd), .A(_82__16_), .Y(Q[16]) );
	BUFX2 BUFX2_26 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .Y(Q[17]) );
	BUFX2 BUFX2_27 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .Y(Q[18]) );
	BUFX2 BUFX2_28 ( .gnd(gnd), .vdd(vdd), .A(_82__19_), .Y(Q[19]) );
	BUFX2 BUFX2_29 ( .gnd(gnd), .vdd(vdd), .A(_82__20_), .Y(Q[20]) );
	BUFX2 BUFX2_30 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .Y(Q[21]) );
	BUFX2 BUFX2_31 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .Y(Q[22]) );
	BUFX2 BUFX2_32 ( .gnd(gnd), .vdd(vdd), .A(_82__23_), .Y(Q[23]) );
	BUFX2 BUFX2_33 ( .gnd(gnd), .vdd(vdd), .A(_82__24_), .Y(Q[24]) );
	BUFX2 BUFX2_34 ( .gnd(gnd), .vdd(vdd), .A(_82__25_), .Y(Q[25]) );
	BUFX2 BUFX2_35 ( .gnd(gnd), .vdd(vdd), .A(_82__26_), .Y(Q[26]) );
	BUFX2 BUFX2_36 ( .gnd(gnd), .vdd(vdd), .A(_82__27_), .Y(Q[27]) );
	BUFX2 BUFX2_37 ( .gnd(gnd), .vdd(vdd), .A(_82__28_), .Y(Q[28]) );
	BUFX2 BUFX2_38 ( .gnd(gnd), .vdd(vdd), .A(_82__29_), .Y(Q[29]) );
	BUFX2 BUFX2_39 ( .gnd(gnd), .vdd(vdd), .A(_82__30_), .Y(Q[30]) );
	BUFX2 BUFX2_40 ( .gnd(gnd), .vdd(vdd), .A(_82__31_), .Y(Q[31]) );
	BUFX2 BUFX2_41 ( .gnd(gnd), .vdd(vdd), .A(_83_), .Y(RCO) );
	DFFPOSX1 DFFPOSX1_19 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_12_), .Q(MODO_reg_7__0_) );
	DFFPOSX1 DFFPOSX1_20 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_14_), .Q(MODO_reg_7__1_) );
	DFFPOSX1 DFFPOSX1_21 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_11_), .Q(MODO_reg_2__0_) );
	DFFPOSX1 DFFPOSX1_22 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_13_), .Q(MODO_reg_2__1_) );
	DFFPOSX1 DFFPOSX1_23 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_3_), .Q(MODO_reg_6__0_) );
	DFFPOSX1 DFFPOSX1_24 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_4_), .Q(MODO_reg_3__1_) );
	DFFPOSX1 DFFPOSX1_25 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_5_), .Q(MODO_reg_7__0_) );
	DFFPOSX1 DFFPOSX1_26 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_6_), .Q(MODO_reg_7__1_) );
	DFFPOSX1 DFFPOSX1_27 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__0_), .Q(MODO_reg_4__0_) );
	DFFPOSX1 DFFPOSX1_28 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_0__1_), .Q(MODO_reg_4__1_) );
	DFFPOSX1 DFFPOSX1_29 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_0__2_), .Q(MODO_reg_6__0_) );
	DFFPOSX1 DFFPOSX1_30 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__3_), .Q(MODO_reg_6__1_) );
	DFFPOSX1 DFFPOSX1_31 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__4_), .Q(MODO_reg_1__0_) );
	DFFPOSX1 DFFPOSX1_32 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__5_), .Q(MODO_reg_1__1_) );
	DFFPOSX1 DFFPOSX1_33 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__6_), .Q(D_reg_0_) );
	DFFPOSX1 DFFPOSX1_34 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__7_), .Q(D_reg_1_) );
	DFFPOSX1 DFFPOSX1_35 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__8_), .Q(D_reg_2_) );
	DFFPOSX1 DFFPOSX1_36 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__9_), .Q(D_reg_3_) );
	DFFPOSX1 DFFPOSX1_37 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_0__10_), .Q(D_reg_4_) );
	DFFPOSX1 DFFPOSX1_38 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_0__11_), .Q(D_reg_5_) );
	DFFPOSX1 DFFPOSX1_39 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__12_), .Q(D_reg_6_) );
	DFFPOSX1 DFFPOSX1_40 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__13_), .Q(D_reg_7_) );
	DFFPOSX1 DFFPOSX1_41 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__14_), .Q(D_reg_8_) );
	DFFPOSX1 DFFPOSX1_42 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__15_), .Q(D_reg_9_) );
	DFFPOSX1 DFFPOSX1_43 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__16_), .Q(D_reg_10_) );
	DFFPOSX1 DFFPOSX1_44 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__17_), .Q(D_reg_11_) );
	DFFPOSX1 DFFPOSX1_45 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__18_), .Q(D_reg_12_) );
	DFFPOSX1 DFFPOSX1_46 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_0__19_), .Q(D_reg_13_) );
	DFFPOSX1 DFFPOSX1_47 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_0__20_), .Q(D_reg_14_) );
	DFFPOSX1 DFFPOSX1_48 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__21_), .Q(D_reg_15_) );
	DFFPOSX1 DFFPOSX1_49 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__22_), .Q(D_reg_16_) );
	DFFPOSX1 DFFPOSX1_50 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_0__23_), .Q(D_reg_17_) );
	DFFPOSX1 DFFPOSX1_51 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_0__24_), .Q(D_reg_18_) );
	DFFPOSX1 DFFPOSX1_52 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_0__25_), .Q(D_reg_25_) );
	DFFPOSX1 DFFPOSX1_53 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_0__26_), .Q(D_reg_26_) );
	DFFPOSX1 DFFPOSX1_54 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_0__27_), .Q(D_reg_27_) );
	DFFPOSX1 DFFPOSX1_55 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_0__28_), .Q(D_reg_28_) );
	DFFPOSX1 DFFPOSX1_56 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_0__29_), .Q(D_reg_29_) );
	DFFPOSX1 DFFPOSX1_57 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_0__30_), .Q(D_reg_30_) );
	DFFPOSX1 DFFPOSX1_58 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_0__31_), .Q(D_reg_31_) );
	DFFPOSX1 DFFPOSX1_59 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_85__0_), .Q(_82__0_) );
	DFFPOSX1 DFFPOSX1_60 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_85__1_), .Q(_82__1_) );
	DFFPOSX1 DFFPOSX1_61 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_85__2_), .Q(_82__2_) );
	DFFPOSX1 DFFPOSX1_62 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_85__3_), .Q(_82__3_) );
	DFFPOSX1 DFFPOSX1_63 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_86_), .Q(cont4b_0_RCO) );
	DFFPOSX1 DFFPOSX1_64 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_84_), .Q(cont4b_0_LOAD) );
	INVX1 INVX1_53 ( .gnd(gnd), .vdd(vdd), .A(_82__7_), .Y(_87_) );
	NAND2X1 NAND2X1_51 ( .gnd(gnd), .vdd(vdd), .A(D_reg_4_), .B(_136_), .Y(_88_) );
	INVX1 INVX1_54 ( .gnd(gnd), .vdd(vdd), .A(_82__6_), .Y(_89_) );
	INVX1 INVX1_55 ( .gnd(gnd), .vdd(vdd), .A(_146_), .Y(_90_) );
	NOR2X1 NOR2X1_21 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_1__0_), .B(_135_), .Y(_91_) );
	INVX1 INVX1_56 ( .gnd(gnd), .vdd(vdd), .A(_82__4_), .Y(_92_) );
	NOR2X1 NOR2X1_22 ( .gnd(gnd), .vdd(vdd), .A(_82__7_), .B(_147_), .Y(_84_) );
	NOR2X1 NOR2X1_23 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_1__0_), .B(MODO_reg_1__1_), .Y(_93_) );
	AOI21X1 AOI21X1_14 ( .gnd(gnd), .vdd(vdd), .A(_120_), .B(_122_), .C(_88_), .Y(_94_) );
	INVX1 INVX1_57 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf3), .Y(_95_) );
	NOR2X1 NOR2X1_24 ( .gnd(gnd), .vdd(vdd), .A(_82__4_), .B(_151_), .Y(_96_) );
	NAND2X1 NAND2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_82__5_), .B(_82__4_), .Y(_97_) );
	NOR2X1 NOR2X1_25 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_180_), .Y(_98_) );
	INVX1 INVX1_58 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_2__0_), .Y(_99_) );
	INVX1 INVX1_59 ( .gnd(gnd), .vdd(vdd), .A(_181_), .Y(_100_) );
	NOR2X1 NOR2X1_26 ( .gnd(gnd), .vdd(vdd), .A(_178_), .B(_182_), .Y(_101_) );
	NAND3X1 NAND3X1_21 ( .gnd(gnd), .vdd(vdd), .A(_82__6_), .B(_82__5_), .C(_82__4_), .Y(_102_) );
	INVX1 INVX1_60 ( .gnd(gnd), .vdd(vdd), .A(_183_), .Y(_103_) );
	NOR2X1 NOR2X1_27 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_2__1_), .B(_179_), .Y(_104_) );
	AND2X2 AND2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_82__7_), .Y(_105_) );
	NAND2X1 NAND2X1_53 ( .gnd(gnd), .vdd(vdd), .A(_158_), .B(_157_), .Y(_106_) );
	NOR2X1 NOR2X1_28 ( .gnd(gnd), .vdd(vdd), .A(_82__9_), .B(_82__8_), .Y(_107_) );
	AOI22X1 AOI22X1_12 ( .gnd(gnd), .vdd(vdd), .A(D_reg_2_), .B(_91_), .C(_93_), .D(_121_), .Y(_108_) );
	AOI21X1 AOI21X1_15 ( .gnd(gnd), .vdd(vdd), .A(_128_), .B(_125_), .C(_88_), .Y(_86_) );
	NAND2X1 NAND2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_162_), .B(_147_), .Y(_109_) );
	INVX1 INVX1_61 ( .gnd(gnd), .vdd(vdd), .A(_82__11_), .Y(_110_) );
	OAI21X1 OAI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_82__2_), .B(_112_), .C(_82__3_), .Y(_111_) );
	AOI21X1 AOI21X1_16 ( .gnd(gnd), .vdd(vdd), .A(_82__5_), .B(_82__4_), .C(_82__6_), .Y(_85__0_) );
	INVX1 INVX1_62 ( .gnd(gnd), .vdd(vdd), .A(_82__10_), .Y(_112_) );
	NOR2X1 NOR2X1_29 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_2__0_), .B(_180_), .Y(_113_) );
	NOR2X1 NOR2X1_30 ( .gnd(gnd), .vdd(vdd), .A(_82__11_), .B(_192_), .Y(_114_) );
	NAND2X1 NAND2X1_55 ( .gnd(gnd), .vdd(vdd), .A(_143_), .B(_171_), .Y(_115_) );
	OR2X2 OR2X2_3 ( .gnd(gnd), .vdd(vdd), .A(_429_), .B(MODO_reg_7__0_), .Y(_116_) );
	AOI22X1 AOI22X1_13 ( .gnd(gnd), .vdd(vdd), .A(_124_), .B(_104_), .C(_100_), .D(_123_), .Y(_117_) );
	AOI21X1 AOI21X1_17 ( .gnd(gnd), .vdd(vdd), .A(_153_), .B(_144_), .C(_133_), .Y(_85__1_) );
	OAI21X1 OAI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_134_), .B(_135_), .C(_155_), .Y(_118_) );
	OAI21X1 OAI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_1__0_), .B(_135_), .C(_163_), .Y(_119_) );
	OAI21X1 OAI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_149_), .B(_163_), .C(_164_), .Y(_120_) );
	NAND3X1 NAND3X1_22 ( .gnd(gnd), .vdd(vdd), .A(_185_), .B(_186_), .C(_187_), .Y(_121_) );
	OAI21X1 OAI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_82__6_), .B(_157_), .C(_82__7_), .Y(_122_) );
	NAND2X1 NAND2X1_56 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_177_), .Y(_123_) );
	AOI22X1 AOI22X1_14 ( .gnd(gnd), .vdd(vdd), .A(D_reg_3_), .B(_91_), .C(_93_), .D(_127_), .Y(_124_) );
	AOI21X1 AOI21X1_18 ( .gnd(gnd), .vdd(vdd), .A(_154_), .B(_156_), .C(_133_), .Y(_85__2_) );
	XOR2X1 XOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_82__3_), .Y(_125_) );
	NAND3X1 NAND3X1_23 ( .gnd(gnd), .vdd(vdd), .A(_82__10_), .B(_82__9_), .C(_82__8_), .Y(_126_) );
	XNOR2X1 XNOR2X1_3 ( .gnd(gnd), .vdd(vdd), .A(_387_), .B(_82__3_), .Y(_127_) );
	AOI22X1 AOI22X1_15 ( .gnd(gnd), .vdd(vdd), .A(_150_), .B(_152_), .C(_145_), .D(_148_), .Y(_128_) );
	NAND2X1 NAND2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_82__10_), .B(_82__9_), .Y(_129_) );
	NAND2X1 NAND2X1_58 ( .gnd(gnd), .vdd(vdd), .A(D_reg_8_), .B(_181_), .Y(_130_) );
	AOI22X1 AOI22X1_16 ( .gnd(gnd), .vdd(vdd), .A(D_reg_5_), .B(_136_), .C(_138_), .D(_159_), .Y(_131_) );
	AOI21X1 AOI21X1_19 ( .gnd(gnd), .vdd(vdd), .A(_160_), .B(_161_), .C(_133_), .Y(_85__3_) );
	DFFPOSX1 DFFPOSX1_65 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_130__0_), .Q(_82__4_) );
	DFFPOSX1 DFFPOSX1_66 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_130__1_), .Q(_82__5_) );
	DFFPOSX1 DFFPOSX1_67 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_130__2_), .Q(_82__6_) );
	DFFPOSX1 DFFPOSX1_68 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_130__3_), .Q(_82__7_) );
	DFFPOSX1 DFFPOSX1_69 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_131_), .Q(cont4b_1_RCO) );
	DFFPOSX1 DFFPOSX1_70 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_129_), .Q(cont4b_1_LOAD) );
	INVX1 INVX1_63 ( .gnd(gnd), .vdd(vdd), .A(_191_), .Y(_135_) );
	NAND2X1 NAND2X1_59 ( .gnd(gnd), .vdd(vdd), .A(_82__9_), .B(_82__8_), .Y(_136_) );
	INVX1 INVX1_64 ( .gnd(gnd), .vdd(vdd), .A(_82__8_), .Y(_137_) );
	INVX1 INVX1_65 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf2), .Y(_138_) );
	NOR2X1 NOR2X1_31 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_2__0_), .B(MODO_reg_2__1_), .Y(_139_) );
	INVX1 INVX1_66 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_3__0_), .Y(_140_) );
	NOR2X1 NOR2X1_32 ( .gnd(gnd), .vdd(vdd), .A(_82__8_), .B(_196_), .Y(_132_) );
	NOR2X1 NOR2X1_33 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .Y(_141_) );
	AOI21X1 AOI21X1_20 ( .gnd(gnd), .vdd(vdd), .A(_165_), .B(_167_), .C(_133_), .Y(_142_) );
	INVX1 INVX1_67 ( .gnd(gnd), .vdd(vdd), .A(_226_), .Y(_143_) );
	NOR2X1 NOR2X1_34 ( .gnd(gnd), .vdd(vdd), .A(_223_), .B(_227_), .Y(_144_) );
	NAND2X1 NAND2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_203_), .B(_202_), .Y(_145_) );
	NOR2X1 NOR2X1_35 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_3__1_), .B(_224_), .Y(_146_) );
	INVX1 INVX1_68 ( .gnd(gnd), .vdd(vdd), .A(_228_), .Y(_147_) );
	INVX1 INVX1_69 ( .gnd(gnd), .vdd(vdd), .A(_82__15_), .Y(_148_) );
	NOR2X1 NOR2X1_36 ( .gnd(gnd), .vdd(vdd), .A(_82__13_), .B(_82__12_), .Y(_149_) );
	NAND3X1 NAND3X1_24 ( .gnd(gnd), .vdd(vdd), .A(_230_), .B(_231_), .C(_232_), .Y(_150_) );
	INVX1 INVX1_70 ( .gnd(gnd), .vdd(vdd), .A(_82__14_), .Y(_151_) );
	NOR2X1 NOR2X1_37 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_3__0_), .B(_225_), .Y(_152_) );
	AND2X2 AND2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_82__11_), .Y(_153_) );
	NAND2X1 NAND2X1_61 ( .gnd(gnd), .vdd(vdd), .A(_207_), .B(_192_), .Y(_154_) );
	NOR2X1 NOR2X1_38 ( .gnd(gnd), .vdd(vdd), .A(_82__15_), .B(_237_), .Y(_155_) );
	AOI22X1 AOI22X1_17 ( .gnd(gnd), .vdd(vdd), .A(D_reg_6_), .B(_136_), .C(_138_), .D(_166_), .Y(_156_) );
	AOI21X1 AOI21X1_21 ( .gnd(gnd), .vdd(vdd), .A(_173_), .B(_170_), .C(_133_), .Y(_134_) );
	NAND2X1 NAND2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_188_), .B(_216_), .Y(_157_) );
	INVX1 INVX1_71 ( .gnd(gnd), .vdd(vdd), .A(_236_), .Y(_158_) );
	OAI21X1 OAI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_179_), .B(_180_), .C(_200_), .Y(_159_) );
	AOI21X1 AOI21X1_22 ( .gnd(gnd), .vdd(vdd), .A(_82__9_), .B(_82__8_), .C(_82__10_), .Y(_133__0_) );
	INVX1 INVX1_72 ( .gnd(gnd), .vdd(vdd), .A(_82__12_), .Y(_160_) );
	NOR2X1 NOR2X1_39 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_3__0_), .B(MODO_reg_3__1_), .Y(_161_) );
	NOR2X1 NOR2X1_40 ( .gnd(gnd), .vdd(vdd), .A(_82__12_), .B(_241_), .Y(_162_) );
	NAND2X1 NAND2X1_63 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_222_), .Y(_163_) );
	OR2X2 OR2X2_4 ( .gnd(gnd), .vdd(vdd), .A(_94_), .B(_98_), .Y(_164_) );
	AOI22X1 AOI22X1_18 ( .gnd(gnd), .vdd(vdd), .A(_169_), .B(_149_), .C(_145_), .D(_168_), .Y(_165_) );
	AOI21X1 AOI21X1_23 ( .gnd(gnd), .vdd(vdd), .A(_198_), .B(_189_), .C(_178_), .Y(_133__1_) );
	OAI21X1 OAI21X1_49 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_2__0_), .B(_180_), .C(_208_), .Y(_166_) );
	OAI21X1 OAI21X1_50 ( .gnd(gnd), .vdd(vdd), .A(_194_), .B(_208_), .C(_209_), .Y(_167_) );
	OAI21X1 OAI21X1_51 ( .gnd(gnd), .vdd(vdd), .A(_82__10_), .B(_202_), .C(_82__11_), .Y(_168_) );
	NAND3X1 NAND3X1_25 ( .gnd(gnd), .vdd(vdd), .A(_82__14_), .B(_82__13_), .C(_82__12_), .Y(_169_) );
	OAI21X1 OAI21X1_52 ( .gnd(gnd), .vdd(vdd), .A(_224_), .B(_225_), .C(_245_), .Y(_170_) );
	NAND2X1 NAND2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_82__14_), .B(_82__13_), .Y(_171_) );
	AOI22X1 AOI22X1_19 ( .gnd(gnd), .vdd(vdd), .A(D_reg_7_), .B(_136_), .C(_138_), .D(_172_), .Y(_172_) );
	AOI21X1 AOI21X1_24 ( .gnd(gnd), .vdd(vdd), .A(_199_), .B(_201_), .C(_178_), .Y(_133__2_) );
	XOR2X1 XOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_142_), .B(_82__7_), .Y(_173_) );
	NAND3X1 NAND3X1_26 ( .gnd(gnd), .vdd(vdd), .A(_275_), .B(_276_), .C(_277_), .Y(_174_) );
	XNOR2X1 XNOR2X1_4 ( .gnd(gnd), .vdd(vdd), .A(_412_), .B(_411_), .Y(_175_) );
	AOI22X1 AOI22X1_20 ( .gnd(gnd), .vdd(vdd), .A(_195_), .B(_197_), .C(_190_), .D(_193_), .Y(_176_) );
	NAND2X1 NAND2X1_65 ( .gnd(gnd), .vdd(vdd), .A(D_reg_12_), .B(_226_), .Y(_177_) );
	NAND2X1 NAND2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_82__13_), .B(_82__12_), .Y(_178_) );
	AOI22X1 AOI22X1_21 ( .gnd(gnd), .vdd(vdd), .A(D_reg_9_), .B(_181_), .C(_183_), .D(_204_), .Y(_179_) );
	AOI21X1 AOI21X1_25 ( .gnd(gnd), .vdd(vdd), .A(_205_), .B(_206_), .C(_178_), .Y(_133__3_) );
	DFFPOSX1 DFFPOSX1_71 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_175__0_), .Q(_82__8_) );
	DFFPOSX1 DFFPOSX1_72 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_175__1_), .Q(_82__9_) );
	DFFPOSX1 DFFPOSX1_73 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_175__2_), .Q(_82__10_) );
	DFFPOSX1 DFFPOSX1_74 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_175__3_), .Q(_82__11_) );
	DFFPOSX1 DFFPOSX1_75 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_176_), .Q(cont4b_2_RCO) );
	DFFPOSX1 DFFPOSX1_76 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_174_), .Q(cont4b_2_LOAD) );
	INVX1 INVX1_73 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf1), .Y(_183_) );
	NAND2X1 NAND2X1_67 ( .gnd(gnd), .vdd(vdd), .A(_248_), .B(_247_), .Y(_184_) );
	INVX1 INVX1_74 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__0_), .Y(_185_) );
	INVX1 INVX1_75 ( .gnd(gnd), .vdd(vdd), .A(_271_), .Y(_186_) );
	NOR2X1 NOR2X1_41 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .Y(_187_) );
	INVX1 INVX1_76 ( .gnd(gnd), .vdd(vdd), .A(_273_), .Y(_188_) );
	NOR2X1 NOR2X1_42 ( .gnd(gnd), .vdd(vdd), .A(_268_), .B(_272_), .Y(_180_) );
	NOR2X1 NOR2X1_43 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__1_), .B(_269_), .Y(_189_) );
	AOI21X1 AOI21X1_26 ( .gnd(gnd), .vdd(vdd), .A(_210_), .B(_212_), .C(_178_), .Y(_190_) );
	INVX1 INVX1_77 ( .gnd(gnd), .vdd(vdd), .A(_82__19_), .Y(_191_) );
	NOR2X1 NOR2X1_44 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .B(_82__16_), .Y(_192_) );
	NAND2X1 NAND2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_252_), .B(_237_), .Y(_193_) );
	NOR2X1 NOR2X1_45 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__0_), .B(_270_), .Y(_194_) );
	INVX1 INVX1_78 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .Y(_195_) );
	INVX1 INVX1_79 ( .gnd(gnd), .vdd(vdd), .A(_281_), .Y(_196_) );
	NOR2X1 NOR2X1_46 ( .gnd(gnd), .vdd(vdd), .A(_82__19_), .B(_282_), .Y(_197_) );
	NAND3X1 NAND3X1_27 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .B(_82__17_), .C(_82__16_), .Y(_198_) );
	INVX1 INVX1_80 ( .gnd(gnd), .vdd(vdd), .A(_82__16_), .Y(_199_) );
	NOR2X1 NOR2X1_47 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__0_), .B(MODO_reg_4__1_), .Y(_200_) );
	AND2X2 AND2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_82__15_), .Y(_201_) );
	NAND2X1 NAND2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_233_), .B(_261_), .Y(_202_) );
	NOR2X1 NOR2X1_48 ( .gnd(gnd), .vdd(vdd), .A(_82__16_), .B(_286_), .Y(_203_) );
	AOI22X1 AOI22X1_22 ( .gnd(gnd), .vdd(vdd), .A(D_reg_10_), .B(_181_), .C(_183_), .D(_211_), .Y(_204_) );
	AOI21X1 AOI21X1_27 ( .gnd(gnd), .vdd(vdd), .A(_218_), .B(_215_), .C(_178_), .Y(_182_) );
	NAND2X1 NAND2X1_70 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_267_), .Y(_205_) );
	INVX1 INVX1_81 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf0), .Y(_206_) );
	OAI21X1 OAI21X1_53 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_3__0_), .B(_225_), .C(_253_), .Y(_207_) );
	AOI21X1 AOI21X1_28 ( .gnd(gnd), .vdd(vdd), .A(_82__13_), .B(_82__12_), .C(_82__14_), .Y(_181__0_) );
	INVX1 INVX1_82 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .Y(_208_) );
	NOR2X1 NOR2X1_49 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .Y(_209_) );
	NOR2X1 NOR2X1_50 ( .gnd(gnd), .vdd(vdd), .A(_313_), .B(_317_), .Y(_210_) );
	NAND2X1 NAND2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .B(_82__17_), .Y(_211_) );
	OR2X2 OR2X2_5 ( .gnd(gnd), .vdd(vdd), .A(_82__1_), .B(_82__0_), .Y(_212_) );
	AOI22X1 AOI22X1_23 ( .gnd(gnd), .vdd(vdd), .A(_214_), .B(_194_), .C(_190_), .D(_213_), .Y(_213_) );
	AOI21X1 AOI21X1_29 ( .gnd(gnd), .vdd(vdd), .A(_243_), .B(_234_), .C(_223_), .Y(_181__1_) );
	OAI21X1 OAI21X1_54 ( .gnd(gnd), .vdd(vdd), .A(_239_), .B(_253_), .C(_254_), .Y(_214_) );
	OAI21X1 OAI21X1_55 ( .gnd(gnd), .vdd(vdd), .A(_82__14_), .B(_247_), .C(_82__15_), .Y(_215_) );
	OAI21X1 OAI21X1_56 ( .gnd(gnd), .vdd(vdd), .A(_269_), .B(_270_), .C(_290_), .Y(_216_) );
	NAND3X1 NAND3X1_28 ( .gnd(gnd), .vdd(vdd), .A(_320_), .B(_321_), .C(_322_), .Y(_217_) );
	OAI21X1 OAI21X1_57 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__0_), .B(_270_), .C(_298_), .Y(_218_) );
	NAND2X1 NAND2X1_72 ( .gnd(gnd), .vdd(vdd), .A(D_reg_16_), .B(_271_), .Y(_219_) );
	AOI22X1 AOI22X1_24 ( .gnd(gnd), .vdd(vdd), .A(D_reg_11_), .B(_181_), .C(_183_), .D(_217_), .Y(_220_) );
	AOI21X1 AOI21X1_30 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_246_), .C(_223_), .Y(_181__2_) );
	XOR2X1 XOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_190_), .B(_82__11_), .Y(_221_) );
	NAND3X1 NAND3X1_29 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .B(_82__21_), .C(_82__20_), .Y(_222_) );
	XNOR2X1 XNOR2X1_5 ( .gnd(gnd), .vdd(vdd), .A(_416_), .B(_410_), .Y(_223_) );
	AOI22X1 AOI22X1_25 ( .gnd(gnd), .vdd(vdd), .A(_240_), .B(_242_), .C(_235_), .D(_238_), .Y(_224_) );
	NAND2X1 NAND2X1_73 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .B(_82__16_), .Y(_225_) );
	NAND2X1 NAND2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_292_), .Y(_226_) );
	AOI22X1 AOI22X1_26 ( .gnd(gnd), .vdd(vdd), .A(D_reg_13_), .B(_226_), .C(_228_), .D(_249_), .Y(_227_) );
	AOI21X1 AOI21X1_31 ( .gnd(gnd), .vdd(vdd), .A(_250_), .B(_251_), .C(_223_), .Y(_181__3_) );
	DFFPOSX1 DFFPOSX1_77 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_220__0_), .Q(_82__12_) );
	DFFPOSX1 DFFPOSX1_78 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_220__1_), .Q(_82__13_) );
	DFFPOSX1 DFFPOSX1_79 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_220__2_), .Q(_82__14_) );
	DFFPOSX1 DFFPOSX1_80 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_220__3_), .Q(_82__15_) );
	DFFPOSX1 DFFPOSX1_81 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_221_), .Q(cont4b_3_RCO) );
	DFFPOSX1 DFFPOSX1_82 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_219_), .Q(cont4b_3_LOAD) );
	INVX1 INVX1_83 ( .gnd(gnd), .vdd(vdd), .A(_316_), .Y(_231_) );
	NAND2X1 NAND2X1_75 ( .gnd(gnd), .vdd(vdd), .A(_297_), .B(_282_), .Y(_232_) );
	INVX1 INVX1_84 ( .gnd(gnd), .vdd(vdd), .A(_318_), .Y(_233_) );
	INVX1 INVX1_85 ( .gnd(gnd), .vdd(vdd), .A(_82__23_), .Y(_234_) );
	NOR2X1 NOR2X1_51 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__1_), .B(_314_), .Y(_235_) );
	INVX1 INVX1_86 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .Y(_236_) );
	NOR2X1 NOR2X1_52 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .B(_82__20_), .Y(_228_) );
	NOR2X1 NOR2X1_53 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .B(_315_), .Y(_237_) );
	AOI21X1 AOI21X1_32 ( .gnd(gnd), .vdd(vdd), .A(_255_), .B(_257_), .C(_223_), .Y(_238_) );
	INVX1 INVX1_87 ( .gnd(gnd), .vdd(vdd), .A(_326_), .Y(_239_) );
	NOR2X1 NOR2X1_54 ( .gnd(gnd), .vdd(vdd), .A(_82__23_), .B(_327_), .Y(_240_) );
	NAND2X1 NAND2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_278_), .B(_306_), .Y(_241_) );
	NOR2X1 NOR2X1_55 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .B(MODO_reg_5__1_), .Y(_242_) );
	INVX1 INVX1_88 ( .gnd(gnd), .vdd(vdd), .A(_82__20_), .Y(_243_) );
	INVX1 INVX1_89 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .Y(_244_) );
	NOR2X1 NOR2X1_56 ( .gnd(gnd), .vdd(vdd), .A(_82__20_), .B(_331_), .Y(_245_) );
	NAND3X1 NAND3X1_30 ( .gnd(gnd), .vdd(vdd), .A(_365_), .B(_366_), .C(_367_), .Y(_368_) );
	INVX1 INVX1_90 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_6__0_), .Y(_247_) );
	NOR2X1 NOR2X1_57 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .Y(_361_) );
	AND2X2 AND2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_82__19_), .Y(_249_) );
	NAND2X1 NAND2X1_77 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_312_), .Y(_250_) );
	NOR2X1 NOR2X1_58 ( .gnd(gnd), .vdd(vdd), .A(_358_), .B(_362_), .Y(_354_) );
	AOI22X1 AOI22X1_27 ( .gnd(gnd), .vdd(vdd), .A(D_reg_14_), .B(_226_), .C(_228_), .D(_256_), .Y(_252_) );
	AOI21X1 AOI21X1_33 ( .gnd(gnd), .vdd(vdd), .A(_263_), .B(_260_), .C(_223_), .Y(_230_) );
	NAND2X1 NAND2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .B(_82__21_), .Y(_253_) );
	INVX1 INVX1_91 ( .gnd(gnd), .vdd(vdd), .A(_361_), .Y(_254_) );
	OAI21X1 OAI21X1_58 ( .gnd(gnd), .vdd(vdd), .A(_284_), .B(_298_), .C(_299_), .Y(_255_) );
	AOI21X1 AOI21X1_34 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .B(_82__16_), .C(_82__18_), .Y(_229__0_) );
	INVX1 INVX1_92 ( .gnd(gnd), .vdd(vdd), .A(_363_), .Y(_256_) );
	NOR2X1 NOR2X1_59 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_6__1_), .B(_359_), .Y(_363_) );
	NOR2X1 NOR2X1_60 ( .gnd(gnd), .vdd(vdd), .A(_82__25_), .B(_82__24_), .Y(_367_) );
	NAND2X1 NAND2X1_79 ( .gnd(gnd), .vdd(vdd), .A(D_reg_20_), .B(_316_), .Y(_259_) );
	OR2X2 OR2X2_6 ( .gnd(gnd), .vdd(vdd), .A(_114_), .B(MODO[0]), .Y(_260_) );
	AOI22X1 AOI22X1_28 ( .gnd(gnd), .vdd(vdd), .A(_259_), .B(_239_), .C(_235_), .D(_258_), .Y(_261_) );
	AOI21X1 AOI21X1_35 ( .gnd(gnd), .vdd(vdd), .A(_288_), .B(_279_), .C(_268_), .Y(_229__1_) );
	OAI21X1 OAI21X1_59 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .B(_292_), .C(_82__19_), .Y(_262_) );
	OAI21X1 OAI21X1_60 ( .gnd(gnd), .vdd(vdd), .A(_314_), .B(_315_), .C(_335_), .Y(_263_) );
	OAI21X1 OAI21X1_61 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .B(_315_), .C(_343_), .Y(_264_) );
	NAND3X1 NAND3X1_31 ( .gnd(gnd), .vdd(vdd), .A(_244_), .B(_256_), .C(_254_), .Y(_265_) );
	OAI21X1 OAI21X1_62 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_343_), .C(_344_), .Y(_266_) );
	NAND2X1 NAND2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .B(_82__20_), .Y(_267_) );
	AOI22X1 AOI22X1_29 ( .gnd(gnd), .vdd(vdd), .A(D_reg_15_), .B(_226_), .C(_228_), .D(_262_), .Y(_268_) );
	AOI21X1 AOI21X1_36 ( .gnd(gnd), .vdd(vdd), .A(_289_), .B(_291_), .C(_268_), .Y(_229__2_) );
	XOR2X1 XOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_238_), .B(_82__15_), .Y(_269_) );
	NAND3X1 NAND3X1_32 ( .gnd(gnd), .vdd(vdd), .A(_82__14_), .B(_82__13_), .C(_82__12_), .Y(_270_) );
	XNOR2X1 XNOR2X1_6 ( .gnd(gnd), .vdd(vdd), .A(_432_), .B(_82__31_), .Y(_271_) );
	AOI22X1 AOI22X1_30 ( .gnd(gnd), .vdd(vdd), .A(_285_), .B(_287_), .C(_280_), .D(_283_), .Y(_272_) );
	NAND2X1 NAND2X1_81 ( .gnd(gnd), .vdd(vdd), .A(_338_), .B(_337_), .Y(_273_) );
	NAND2X1 NAND2X1_82 ( .gnd(gnd), .vdd(vdd), .A(_342_), .B(_327_), .Y(_274_) );
	AOI22X1 AOI22X1_31 ( .gnd(gnd), .vdd(vdd), .A(D_reg_17_), .B(_271_), .C(_273_), .D(_294_), .Y(_275_) );
	AOI21X1 AOI21X1_37 ( .gnd(gnd), .vdd(vdd), .A(_295_), .B(_296_), .C(_268_), .Y(_229__3_) );
	DFFPOSX1 DFFPOSX1_83 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_265__0_), .Q(_82__16_) );
	DFFPOSX1 DFFPOSX1_84 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_265__1_), .Q(_82__17_) );
	DFFPOSX1 DFFPOSX1_85 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_265__2_), .Q(_82__18_) );
	DFFPOSX1 DFFPOSX1_86 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf4), .D(_265__3_), .Q(_82__19_) );
	DFFPOSX1 DFFPOSX1_87 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf3), .D(_266_), .Q(cont4b_4_RCO) );
	DFFPOSX1 DFFPOSX1_88 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf2), .D(_264_), .Q(cont4b_4_LOAD) );
	INVX1 INVX1_93 ( .gnd(gnd), .vdd(vdd), .A(_82__27_), .Y(_365_) );
	NAND2X1 NAND2X1_83 ( .gnd(gnd), .vdd(vdd), .A(_323_), .B(_351_), .Y(_280_) );
	INVX1 INVX1_94 ( .gnd(gnd), .vdd(vdd), .A(_82__26_), .Y(_366_) );
	INVX1 INVX1_95 ( .gnd(gnd), .vdd(vdd), .A(_371_), .Y(_372_) );
	NOR2X1 NOR2X1_61 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_6__0_), .B(_360_), .Y(_370_) );
	INVX1 INVX1_96 ( .gnd(gnd), .vdd(vdd), .A(_82__24_), .Y(_284_) );
	NOR2X1 NOR2X1_62 ( .gnd(gnd), .vdd(vdd), .A(_82__27_), .B(_372_), .Y(_276_) );
	NOR2X1 NOR2X1_63 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_6__0_), .B(MODO_reg_6__1_), .Y(_374_) );
	AOI21X1 AOI21X1_38 ( .gnd(gnd), .vdd(vdd), .A(_300_), .B(_302_), .C(_268_), .Y(_286_) );
	INVX1 INVX1_97 ( .gnd(gnd), .vdd(vdd), .A(_286_), .Y(_287_) );
	NOR2X1 NOR2X1_64 ( .gnd(gnd), .vdd(vdd), .A(_82__24_), .B(_376_), .Y(_288_) );
	NAND2X1 NAND2X1_84 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_357_), .Y(_358_) );
	NOR2X1 NOR2X1_65 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__1_), .B(_281_), .Y(_290_) );
	INVX1 INVX1_98 ( .gnd(gnd), .vdd(vdd), .A(_82__19_), .Y(_291_) );
	INVX1 INVX1_99 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .Y(_292_) );
	NOR2X1 NOR2X1_66 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .B(_82__16_), .Y(_293_) );
	NAND3X1 NAND3X1_33 ( .gnd(gnd), .vdd(vdd), .A(_291_), .B(_292_), .C(_293_), .Y(_294_) );
	INVX1 INVX1_100 ( .gnd(gnd), .vdd(vdd), .A(_294_), .Y(_295_) );
	NOR2X1 NOR2X1_67 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__0_), .B(MODO_reg_4__1_), .Y(_296_) );
	AND2X2 AND2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_82__23_), .Y(_297_) );
	NAND2X1 NAND2X1_85 ( .gnd(gnd), .vdd(vdd), .A(_82__26_), .B(_82__25_), .Y(_298_) );
	NOR2X1 NOR2X1_68 ( .gnd(gnd), .vdd(vdd), .A(_82__16_), .B(_298_), .Y(_299_) );
	AOI22X1 AOI22X1_32 ( .gnd(gnd), .vdd(vdd), .A(D_reg_18_), .B(_271_), .C(_273_), .D(_301_), .Y(_300_) );
	AOI21X1 AOI21X1_39 ( .gnd(gnd), .vdd(vdd), .A(_308_), .B(_305_), .C(_268_), .Y(_278_) );
	NAND2X1 NAND2X1_86 ( .gnd(gnd), .vdd(vdd), .A(D_reg_24_), .B(_361_), .Y(_301_) );
	INVX1 INVX1_101 ( .gnd(gnd), .vdd(vdd), .A(_82__16_), .Y(_302_) );
	OAI21X1 OAI21X1_63 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .B(_337_), .C(_82__23_), .Y(_303_) );
	AOI21X1 AOI21X1_40 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .B(_82__20_), .C(_82__22_), .Y(_277__0_) );
	INVX1 INVX1_102 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .Y(_304_) );
	NOR2X1 NOR2X1_69 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_302_), .Y(_305_) );
	NOR2X1 NOR2X1_70 ( .gnd(gnd), .vdd(vdd), .A(_293_), .B(_305_), .Y(_306_) );
	NAND2X1 NAND2X1_87 ( .gnd(gnd), .vdd(vdd), .A(_82__25_), .B(_82__24_), .Y(_307_) );
	OR2X2 OR2X2_7 ( .gnd(gnd), .vdd(vdd), .A(_139_), .B(_143_), .Y(_308_) );
	AOI22X1 AOI22X1_33 ( .gnd(gnd), .vdd(vdd), .A(_304_), .B(_284_), .C(_280_), .D(_303_), .Y(_309_) );
	AOI21X1 AOI21X1_41 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_324_), .C(_313_), .Y(_277__1_) );
	OAI21X1 OAI21X1_64 ( .gnd(gnd), .vdd(vdd), .A(_359_), .B(_360_), .C(_380_), .Y(_310_) );
	OAI21X1 OAI21X1_65 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_4__0_), .B(_282_), .C(_310_), .Y(_311_) );
	OAI21X1 OAI21X1_66 ( .gnd(gnd), .vdd(vdd), .A(_296_), .B(_310_), .C(_311_), .Y(_312_) );
	NAND3X1 NAND3X1_34 ( .gnd(gnd), .vdd(vdd), .A(_292_), .B(_304_), .C(_302_), .Y(_313_) );
	OAI21X1 OAI21X1_67 ( .gnd(gnd), .vdd(vdd), .A(_82__17_), .B(_82__16_), .C(_82__18_), .Y(_314_) );
	NAND2X1 NAND2X1_88 ( .gnd(gnd), .vdd(vdd), .A(_383_), .B(_382_), .Y(_384_) );
	AOI22X1 AOI22X1_34 ( .gnd(gnd), .vdd(vdd), .A(D_reg_19_), .B(_271_), .C(_273_), .D(_307_), .Y(_316_) );
	AOI21X1 AOI21X1_42 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_336_), .C(_313_), .Y(_277__2_) );
	XOR2X1 XOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_286_), .B(_82__19_), .Y(_317_) );
	NAND3X1 NAND3X1_35 ( .gnd(gnd), .vdd(vdd), .A(_82__18_), .B(_82__17_), .C(_82__16_), .Y(_318_) );
	XNOR2X1 XNOR2X1_7 ( .gnd(gnd), .vdd(vdd), .A(_97_), .B(_96_), .Y(_319_) );
	AOI22X1 AOI22X1_35 ( .gnd(gnd), .vdd(vdd), .A(_330_), .B(_332_), .C(_325_), .D(_328_), .Y(_320_) );
	NAND2X1 NAND2X1_89 ( .gnd(gnd), .vdd(vdd), .A(_82__19_), .B(_313_), .Y(_321_) );
	NAND2X1 NAND2X1_90 ( .gnd(gnd), .vdd(vdd), .A(_294_), .B(_321_), .Y(_322_) );
	AOI22X1 AOI22X1_36 ( .gnd(gnd), .vdd(vdd), .A(D_reg_21_), .B(_316_), .C(_318_), .D(_339_), .Y(_323_) );
	AOI21X1 AOI21X1_43 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_341_), .C(_313_), .Y(_277__3_) );
	DFFPOSX1 DFFPOSX1_89 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf1), .D(_310__0_), .Q(_82__20_) );
	DFFPOSX1 DFFPOSX1_90 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf0), .D(_310__1_), .Q(_82__21_) );
	DFFPOSX1 DFFPOSX1_91 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf8), .D(_310__2_), .Q(_82__22_) );
	DFFPOSX1 DFFPOSX1_92 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf7), .D(_310__3_), .Q(_82__23_) );
	DFFPOSX1 DFFPOSX1_93 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf6), .D(_311_), .Q(cont4b_5_RCO) );
	DFFPOSX1 DFFPOSX1_94 ( .gnd(gnd), .vdd(vdd), .CLK(clk_bF_buf5), .D(_309_), .Q(cont4b_5_LOAD) );
	INVX1 INVX1_103 ( .gnd(gnd), .vdd(vdd), .A(RESET_bF_buf7), .Y(_327_) );
	NAND2X1 NAND2X1_91 ( .gnd(gnd), .vdd(vdd), .A(ENABLE), .B(_327_), .Y(_328_) );
	INVX1 INVX1_104 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .Y(_329_) );
	INVX1 INVX1_105 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__1_), .Y(_330_) );
	NOR2X1 NOR2X1_71 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .Y(_331_) );
	INVX1 INVX1_106 ( .gnd(gnd), .vdd(vdd), .A(_331_), .Y(_332_) );
	NOR2X1 NOR2X1_72 ( .gnd(gnd), .vdd(vdd), .A(_328_), .B(_332_), .Y(_324_) );
	NOR2X1 NOR2X1_73 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .B(_330_), .Y(_333_) );
	AOI21X1 AOI21X1_44 ( .gnd(gnd), .vdd(vdd), .A(_345_), .B(_347_), .C(_313_), .Y(_334_) );
	INVX1 INVX1_107 ( .gnd(gnd), .vdd(vdd), .A(_334_), .Y(_335_) );
	NOR2X1 NOR2X1_74 ( .gnd(gnd), .vdd(vdd), .A(_82__23_), .B(_335_), .Y(_336_) );
	NAND2X1 NAND2X1_92 ( .gnd(gnd), .vdd(vdd), .A(_333_), .B(_336_), .Y(_337_) );
	NOR2X1 NOR2X1_75 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__1_), .B(_329_), .Y(_338_) );
	INVX1 INVX1_108 ( .gnd(gnd), .vdd(vdd), .A(_82__23_), .Y(_339_) );
	INVX1 INVX1_109 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .Y(_340_) );
	NOR2X1 NOR2X1_76 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .B(_82__20_), .Y(_341_) );
	NAND3X1 NAND3X1_36 ( .gnd(gnd), .vdd(vdd), .A(_339_), .B(_340_), .C(_341_), .Y(_342_) );
	INVX1 INVX1_110 ( .gnd(gnd), .vdd(vdd), .A(_342_), .Y(_343_) );
	NOR2X1 NOR2X1_77 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .B(MODO_reg_5__1_), .Y(_344_) );
	AND2X2 AND2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_374_), .B(_82__27_), .Y(_345_) );
	NAND2X1 NAND2X1_93 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .B(_82__21_), .Y(_346_) );
	NOR2X1 NOR2X1_78 ( .gnd(gnd), .vdd(vdd), .A(_82__20_), .B(_346_), .Y(_347_) );
	AOI22X1 AOI22X1_37 ( .gnd(gnd), .vdd(vdd), .A(D_reg_22_), .B(_316_), .C(_318_), .D(_346_), .Y(_348_) );
	AOI21X1 AOI21X1_45 ( .gnd(gnd), .vdd(vdd), .A(_353_), .B(_350_), .C(_313_), .Y(_326_) );
	NAND2X1 NAND2X1_94 ( .gnd(gnd), .vdd(vdd), .A(D_reg_20_), .B(_331_), .Y(_349_) );
	INVX1 INVX1_111 ( .gnd(gnd), .vdd(vdd), .A(_82__20_), .Y(_350_) );
	OAI21X1 OAI21X1_68 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_330_), .C(_350_), .Y(_351_) );
	AOI21X1 AOI21X1_46 ( .gnd(gnd), .vdd(vdd), .A(_82__25_), .B(_82__24_), .C(_82__26_), .Y(_371_) );
	INVX1 INVX1_112 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .Y(_352_) );
	NOR2X1 NOR2X1_79 ( .gnd(gnd), .vdd(vdd), .A(_352_), .B(_350_), .Y(_353_) );
	NOR2X1 NOR2X1_80 ( .gnd(gnd), .vdd(vdd), .A(_341_), .B(_353_), .Y(_354_) );
	NAND2X1 NAND2X1_95 ( .gnd(gnd), .vdd(vdd), .A(_329_), .B(_354_), .Y(_355_) );
	OR2X2 OR2X2_8 ( .gnd(gnd), .vdd(vdd), .A(_82__5_), .B(_82__4_), .Y(_356_) );
	AOI22X1 AOI22X1_38 ( .gnd(gnd), .vdd(vdd), .A(_349_), .B(_329_), .C(_325_), .D(_348_), .Y(_357_) );
	AOI21X1 AOI21X1_47 ( .gnd(gnd), .vdd(vdd), .A(_378_), .B(_369_), .C(_358_), .Y(_356_) );
	OAI21X1 OAI21X1_69 ( .gnd(gnd), .vdd(vdd), .A(_350_), .B(_346_), .C(_335_), .Y(_358_) );
	OAI21X1 OAI21X1_70 ( .gnd(gnd), .vdd(vdd), .A(MODO_reg_5__0_), .B(_330_), .C(_358_), .Y(_359_) );
	OAI21X1 OAI21X1_71 ( .gnd(gnd), .vdd(vdd), .A(_344_), .B(_358_), .C(_359_), .Y(_360_) );
	NAND3X1 NAND3X1_37 ( .gnd(gnd), .vdd(vdd), .A(_340_), .B(_352_), .C(_350_), .Y(_361_) );
	OAI21X1 OAI21X1_72 ( .gnd(gnd), .vdd(vdd), .A(_82__21_), .B(_82__20_), .C(_82__22_), .Y(_362_) );
	NAND2X1 NAND2X1_96 ( .gnd(gnd), .vdd(vdd), .A(_362_), .B(_361_), .Y(_363_) );
	AOI22X1 AOI22X1_39 ( .gnd(gnd), .vdd(vdd), .A(D_reg_23_), .B(_316_), .C(_318_), .D(_352_), .Y(_364_) );
	AOI21X1 AOI21X1_48 ( .gnd(gnd), .vdd(vdd), .A(_379_), .B(_381_), .C(_358_), .Y(_355__0_) );
	XOR2X1 XOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_334_), .B(_82__23_), .Y(_365_) );
	NAND3X1 NAND3X1_38 ( .gnd(gnd), .vdd(vdd), .A(_82__22_), .B(_82__21_), .C(_82__20_), .Y(_366_) );
	XNOR2X1 XNOR2X1_8 ( .gnd(gnd), .vdd(vdd), .A(_101_), .B(_95_), .Y(_367_) );
	AOI22X1 AOI22X1_40 ( .gnd(gnd), .vdd(vdd), .A(_375_), .B(_377_), .C(_370_), .D(_373_), .Y(_368_) );
endmodule
