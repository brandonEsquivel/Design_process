*** SPICE deck for cell NAND3{lay} from library gates
*** Created on lun dic 07, 2020 00:24:56
*** Last revised on mar dic 08, 2020 16:13:20
*** Written on mar dic 08, 2020 16:13:30 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** TOP LEVEL CELL: NAND3{lay}
Mnmos@4 net@17 A gnd gnd N L=0.4U W=1U AS=6.02P AD=0.78P PS=17.4U PD=3.2U
Mnmos@5 net@16 B net@17 gnd N L=0.4U W=1U AS=0.78P AD=0.78P PS=3.2U PD=3.2U
Mnmos@6 Y_NAND3 C net@16 gnd N L=0.4U W=1U AS=0.78P AD=2.12P PS=3.2U PD=6.1U
Mpmos@3 Y_NAND3 A vdd vdd P L=0.4U W=2U AS=8.793P AD=2.12P PS=13.533U PD=6.1U
Mpmos@4 vdd B Y_NAND3 vdd P L=0.4U W=2U AS=2.12P AD=8.793P PS=6.1U PD=13.533U
Mpmos@5 Y_NAND3 C vdd vdd P L=0.4U W=2U AS=8.793P AD=2.12P PS=13.533U PD=6.1U

* Spice Code nodes in cell cell 'NAND3{lay}'
vdd VDD 0 DC 5
vin A 0 pulse(0 5 10n 0.5n 0.5n 20n)
vin2 B 0 pulse(0 5 30n 0.5n 0.5n 50n)
vin3 C 0 pulse(0 5 40n 0.5n 0.5n 60n)
.TRAN 0 80n
.MODEL N NMOS
.MODEL P PMOS
.end
.END
